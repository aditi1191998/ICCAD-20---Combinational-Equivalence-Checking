module top(\A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,
        \A[0][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,
        \A[1][0] ,\A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,
        \A[2][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,
        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ,\O[19] ,
        \O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,\O[10] ,\O[9] ,
        \O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,\O[0] );
input \A[0][9] ,\A[0][8] ,\A[0][7] ,\A[0][6] ,\A[0][5] ,\A[0][4] ,\A[0][3] ,\A[0][2] ,\A[0][1] ,
        \A[0][0] ,\A[1][9] ,\A[1][8] ,\A[1][7] ,\A[1][6] ,\A[1][5] ,\A[1][4] ,\A[1][3] ,\A[1][2] ,\A[1][1] ,
        \A[1][0] ,\A[2][9] ,\A[2][8] ,\A[2][7] ,\A[2][6] ,\A[2][5] ,\A[2][4] ,\A[2][3] ,\A[2][2] ,\A[2][1] ,
        \A[2][0] ,\B[9] ,\B[8] ,\B[7] ,\B[6] ,\B[5] ,\B[4] ,\B[3] ,\B[2] ,\B[1] ,
        \B[0] ,\I[7] ,\I[6] ,\I[5] ,\I[4] ,\I[3] ,\I[2] ,\I[1] ,\I[0] ;
output \O[19] ,\O[18] ,\O[17] ,\O[16] ,\O[15] ,\O[14] ,\O[13] ,\O[12] ,\O[11] ,
        \O[10] ,\O[9] ,\O[8] ,\O[7] ,\O[6] ,\O[5] ,\O[4] ,\O[3] ,\O[2] ,\O[1] ,
        \O[0] ;

wire \69_ZERO , \70_ONE , \71 , \72 , \73 , \74 , \75 , \76 , \77 ,
         \78 , \79 , \80 , \81 , \82 , \83 , \84 , \85 , \86 , \87 ,
         \88 , \89 , \90 , \91 , \92 , \93 , \94 , \95 , \96 , \97 ,
         \98 , \99 , \100 , \101 , \102 , \103 , \104 , \105 , \106 , \107 ,
         \108 , \109 , \110 , \111 , \112 , \113 , \114 , \115 , \116 , \117 ,
         \118 , \119 , \120 , \121 , \122 , \123 , \124 , \125 , \126 , \127 ,
         \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 , \136 , \137 ,
         \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 , \146 , \147 ,
         \148 , \149 , \150 , \151 , \152 , \153 , \154 , \155 , \156 , \157 ,
         \158 , \159 , \160 , \161 , \162 , \163 , \164 , \165 , \166 , \167 ,
         \168 , \169 , \170 , \171 , \172 , \173 , \174 , \175 , \176 , \177 ,
         \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 , \186 , \187 ,
         \188 , \189 , \190 , \191 , \192 , \193 , \194 , \195 , \196 , \197 ,
         \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 , \206 , \207 ,
         \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 , \216 , \217 ,
         \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 , \226 , \227 ,
         \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 , \236 , \237 ,
         \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 , \246 , \247 ,
         \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 , \256 , \257 ,
         \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 , \266 , \267 ,
         \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 , \276 , \277 ,
         \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 , \286 , \287 ,
         \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 , \296 , \297 ,
         \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 , \306 , \307 ,
         \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 , \316 , \317 ,
         \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 , \326 , \327 ,
         \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 , \336 , \337 ,
         \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 , \346 , \347 ,
         \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 , \356 , \357 ,
         \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 , \366 , \367 ,
         \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 , \376 , \377 ,
         \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 , \386 , \387 ,
         \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 , \396 , \397 ,
         \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 , \406 , \407 ,
         \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 , \416 , \417 ,
         \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 , \426 , \427 ,
         \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 , \436 , \437 ,
         \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 , \446 , \447 ,
         \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 , \456 , \457 ,
         \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 , \466 , \467 ,
         \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 , \476 , \477 ,
         \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 , \486 , \487 ,
         \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 , \496 , \497 ,
         \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 , \506 , \507 ,
         \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 , \516 , \517 ,
         \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 , \526 , \527 ,
         \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 , \536 , \537 ,
         \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 , \546 , \547 ,
         \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 , \556 , \557 ,
         \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 , \566 , \567 ,
         \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 , \576 , \577 ,
         \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 , \586 , \587 ,
         \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 , \596 , \597 ,
         \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 , \606 , \607 ,
         \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 , \616 , \617 ,
         \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 , \626 , \627 ,
         \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 , \636 , \637 ,
         \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 , \646 , \647 ,
         \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,
         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,
         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 ;
buf \U$labaj121 ( \O[19] , \934 );
buf \U$labaj122 ( \O[18] , \940 );
buf \U$labaj123 ( \O[17] , \960 );
buf \U$labaj124 ( \O[16] , \1067 );
buf \U$labaj125 ( \O[15] , \979 );
buf \U$labaj126 ( \O[14] , \1068 );
buf \U$labaj127 ( \O[13] , \991 );
buf \U$labaj128 ( \O[12] , \1069 );
buf \U$labaj129 ( \O[11] , \1004 );
buf \U$labaj130 ( \O[10] , \1011 );
buf \U$labaj131 ( \O[9] , \1018 );
buf \U$labaj132 ( \O[8] , \1024 );
buf \U$labaj133 ( \O[7] , \1033 );
buf \U$labaj134 ( \O[6] , \1041 );
buf \U$labaj135 ( \O[5] , \1047 );
buf \U$labaj136 ( \O[4] , \1053 );
buf \U$labaj137 ( \O[3] , \1059 );
buf \U$labaj138 ( \O[2] , \1061 );
buf \U$labaj139 ( \O[1] , \1065 );
buf \U$labaj140 ( \O[0] , \1066 );
nor \g11962/U$1 ( \71 , \I[1] , \I[0] );
not \g12001/U$3 ( \72 , \71 );
not \g12001/U$4 ( \73 , \A[0][9] );
or \g12001/U$2 ( \74 , \72 , \73 );
and \g710/U$2 ( \75 , \A[1][9] , \I[0] );
and \g710/U$3 ( \76 , \A[2][9] , \I[1] );
nor \g710/U$1 ( \77 , \75 , \76 );
nand \g12001/U$1 ( \78 , \74 , \77 );
buf \g674/U$1 ( \79 , \78 );
not \g11989/U$2 ( \80 , \A[0][7] );
nor \g11989/U$1 ( \81 , \80 , \I[0] , \I[1] );
nand \g723/U$1 ( \82 , \A[2][7] , \I[1] );
nand \g724/U$1 ( \83 , \A[1][7] , \I[0] );
nand \g709/U$1 ( \84 , \82 , \83 );
nor \g677/U$1 ( \85 , \81 , \84 );
not \g676/U$1 ( \86 , \85 );
not \g11877/U$3 ( \87 , \A[0][5] );
nor \g3/U$1 ( \88 , \I[1] , \I[0] );
not \g11877/U$4 ( \89 , \88 );
or \g11877/U$2 ( \90 , \87 , \89 );
and \g707/U$2 ( \91 , \A[1][5] , \I[0] );
and \g707/U$3 ( \92 , \A[2][5] , \I[1] );
nor \g707/U$1 ( \93 , \91 , \92 );
nand \g11877/U$1 ( \94 , \90 , \93 );
buf \g678/U$1 ( \95 , \94 );
nor \g11960/U$1 ( \96 , \I[1] , \I[0] );
not \g12002/U$3 ( \97 , \96 );
not \g12002/U$4 ( \98 , \A[0][2] );
or \g12002/U$2 ( \99 , \97 , \98 );
and \g704/U$2 ( \100 , \A[1][2] , \I[0] );
and \g704/U$3 ( \101 , \A[2][2] , \I[1] );
nor \g704/U$1 ( \102 , \100 , \101 );
nand \g12002/U$1 ( \103 , \99 , \102 );
buf \g680/U$1 ( \104 , \103 );
not \g11939/U$2 ( \105 , \A[0][1] );
nor \g11939/U$1 ( \106 , \105 , \I[0] , \I[1] );
nand \g718/U$1 ( \107 , \A[2][1] , \I[1] );
nand \g720/U$1 ( \108 , \A[1][1] , \I[0] );
nand \g706/U$1 ( \109 , \107 , \108 );
nor \g683/U$1 ( \110 , \106 , \109 );
not \g682/U$1 ( \111 , \110 );
nor \g11964/U$1 ( \112 , \I[1] , \I[0] );
nand \g11963/U$1 ( \113 , \112 , \A[0][0] );
and \g708/U$2 ( \114 , \A[1][0] , \I[0] );
and \g708/U$3 ( \115 , \A[2][0] , \I[1] );
nor \g708/U$1 ( \116 , \114 , \115 );
nand \g685/U$1 ( \117 , \113 , \116 );
buf \g684/U$1 ( \118 , \117 );
nor \g11968/U$1 ( \119 , \I[1] , \I[0] );
not \g12005/U$3 ( \120 , \119 );
not \g12005/U$4 ( \121 , \A[0][4] );
or \g12005/U$2 ( \122 , \120 , \121 );
and \g711/U$2 ( \123 , \A[1][4] , \I[0] );
and \g711/U$3 ( \124 , \A[2][4] , \I[1] );
nor \g711/U$1 ( \125 , \123 , \124 );
nand \g12005/U$1 ( \126 , \122 , \125 );
buf \g687/U$1 ( \127 , \126 );
nor \g11970/U$1 ( \128 , \I[1] , \I[0] );
not \g12006/U$3 ( \129 , \128 );
not \g12006/U$4 ( \130 , \A[0][6] );
or \g12006/U$2 ( \131 , \129 , \130 );
and \g703/U$2 ( \132 , \A[1][6] , \I[0] );
and \g703/U$3 ( \133 , \A[2][6] , \I[1] );
nor \g703/U$1 ( \134 , \132 , \133 );
nand \g12006/U$1 ( \135 , \131 , \134 );
buf \g689/U$1 ( \136 , \135 );
not \g735/U$1 ( \137 , \A[0][3] );
nor \g701/U$1 ( \138 , \137 , \I[0] , \I[1] );
nand \g715/U$1 ( \139 , \A[2][3] , \I[1] );
nand \g714/U$1 ( \140 , \A[1][3] , \I[0] );
nand \g712/U$1 ( \141 , \139 , \140 );
nor \g692/U$1 ( \142 , \138 , \141 );
not \g691/U$1 ( \143 , \142 );
and \g705/U$2 ( \144 , \A[1][8] , \I[0] );
and \g705/U$3 ( \145 , \A[2][8] , \I[1] );
nor \g705/U$1 ( \146 , \144 , \145 );
nand \mul_6_19_g11706/U$1 ( \147 , \79 , \B[8] );
nor \g11966/U$1 ( \148 , \I[1] , \I[0] );
not \g12004/U$3 ( \149 , \148 );
not \g12004/U$4 ( \150 , \A[0][8] );
or \g12004/U$2 ( \151 , \149 , \150 );
nand \g12004/U$1 ( \152 , \151 , \146 );
buf \mul_6_19_g11756/U$1 ( \153 , \152 );
nand \mul_6_19_g11621/U$1 ( \154 , \153 , \B[9] );
xor \mul_6_19_g11476/U$4 ( \155 , \147 , \154 );
nand \mul_6_19_g11687/U$1 ( \156 , \79 , \B[7] );
nand \mul_6_19_g11634/U$1 ( \157 , \86 , \B[9] );
xor \mul_6_19_g11520/U$4 ( \158 , \156 , \157 );
nand \mul_6_19_g11667/U$1 ( \159 , \153 , \B[8] );
and \mul_6_19_g11520/U$3 ( \160 , \158 , \159 );
and \mul_6_19_g11520/U$5 ( \161 , \156 , \157 );
or \mul_6_19_g11520/U$2 ( \162 , \160 , \161 );
and \mul_6_19_g11476/U$3 ( \163 , \155 , \162 );
and \mul_6_19_g11476/U$5 ( \164 , \147 , \154 );
or \mul_6_19_g11476/U$2 ( \165 , \163 , \164 );
nand \mul_6_19_g11753/U$1 ( \166 , \79 , \B[9] );
nand \mul_6_19_g11454/U$1 ( \167 , \165 , \166 );
not \mul_6_19_g11245/U$3 ( \168 , \167 );
nand \mul_6_19_g11660/U$1 ( \169 , \95 , \B[7] );
nand \mul_6_19_g11676/U$1 ( \170 , \127 , \B[8] );
xor \mul_6_19_g11986/U$1 ( \171 , \169 , \170 );
nand \mul_6_19_g11630/U$1 ( \172 , \86 , \B[5] );
xor \mul_6_19_g11986/U$1_r1 ( \173 , \171 , \172 );
nand \mul_6_19_g11985/U$1 ( \174 , \79 , \B[3] );
nand \mul_6_19_g11715/U$1 ( \175 , \152 , \B[4] );
xor \g11956/U$1 ( \176 , \174 , \175 );
and \mul_6_19_g11689/U$1 ( \177 , \136 , \B[6] );
xnor \g11956/U$1_r1 ( \178 , \176 , \177 );
and \mul_6_19_g11456/U$2 ( \179 , \173 , \178 );
nand \mul_6_19_g11662/U$1 ( \180 , \143 , \B[8] );
nand \mul_6_19_g11869/U$1 ( \181 , \127 , \B[7] );
xor \mul_6_19_g11519/U$4 ( \182 , \180 , \181 );
and \mul_6_19_g11703/U$1 ( \183 , \79 , \B[1] );
and \mul_6_19_g11718/U$1 ( \184 , \152 , \B[2] );
nand \mul_6_19_g11610/U$1 ( \185 , \183 , \184 );
and \mul_6_19_g11519/U$3 ( \186 , \182 , \185 );
and \mul_6_19_g11519/U$5 ( \187 , \180 , \181 );
or \mul_6_19_g11519/U$2 ( \188 , \186 , \187 );
nor \mul_6_19_g11456/U$1 ( \189 , \179 , \188 );
not \fopt11893/U$1 ( \190 , \178 );
not \mul_6_19_g11529/U$1 ( \191 , \173 );
and \mul_6_19_g11475/U$2 ( \192 , \190 , \191 );
nor \mul_6_19_g11433/U$1 ( \193 , \189 , \192 );
not \mul_6_19_g11340/U$3 ( \194 , \193 );
nand \mul_6_19_g11709/U$1 ( \195 , \95 , \B[8] );
nand \mul_6_19_g11868/U$1 ( \196 , \127 , \B[9] );
xor \mul_6_19_g11512/U$1 ( \197 , \195 , \196 );
nand \mul_6_19_g11742/U$1 ( \198 , \86 , \B[6] );
xor \mul_6_19_g11512/U$1_r1 ( \199 , \197 , \198 );
buf \mul_6_19_g11754/U$1 ( \200 , \143 );
nand \mul_6_19_g11727/U$1 ( \201 , \200 , \B[9] );
nand \mul_6_19_g11674/U$1 ( \202 , \152 , \B[3] );
nand \mul_6_19_g11935/U$1 ( \203 , \136 , \B[5] );
xor \mul_6_19_g11510/U$4 ( \204 , \202 , \203 );
nand \mul_6_19_g11701/U$1 ( \205 , \79 , \B[2] );
and \mul_6_19_g11510/U$3 ( \206 , \204 , \205 );
and \mul_6_19_g11510/U$5 ( \207 , \202 , \203 );
or \mul_6_19_g11510/U$2 ( \208 , \206 , \207 );
xor \mul_6_19_g11439/U$4 ( \209 , \201 , \208 );
nand \mul_6_19_g11635/U$1 ( \210 , \95 , \B[6] );
nand \mul_6_19_g11744/U$1 ( \211 , \104 , \B[9] );
xor \mul_6_19_g11532/U$4 ( \212 , \210 , \211 );
nand \mul_6_19_g11751/U$1 ( \213 , \86 , \B[4] );
and \mul_6_19_g11532/U$3 ( \214 , \212 , \213 );
and \mul_6_19_g11532/U$5 ( \215 , \210 , \211 );
or \mul_6_19_g11532/U$2 ( \216 , \214 , \215 );
and \mul_6_19_g11439/U$3 ( \217 , \209 , \216 );
and \mul_6_19_g11439/U$5 ( \218 , \201 , \208 );
or \mul_6_19_g11439/U$2 ( \219 , \217 , \218 );
xor \mul_6_19_g11402/U$1 ( \220 , \199 , \219 );
not \mul_6_19_g11561/U$3 ( \221 , \175 );
not \mul_6_19_g11561/U$4 ( \222 , \174 );
or \mul_6_19_g11561/U$2 ( \223 , \221 , \222 );
nand \mul_6_19_g11561/U$1 ( \224 , \223 , \177 );
not \mul_6_19_g11602/U$2 ( \225 , \174 );
not \mul_6_19_g11714/U$1 ( \226 , \175 );
nand \mul_6_19_g11602/U$1 ( \227 , \225 , \226 );
nand \mul_6_19_g11533/U$1 ( \228 , \224 , \227 );
not \mul_6_19_g11526/U$1 ( \229 , \228 );
not \mul_6_19_g11492/U$3 ( \230 , \229 );
and \g11982/U$1 ( \231 , \169 , \172 );
or \g11981/U$2 ( \232 , \231 , \170 );
or \mul_6_19_g11784/U$1 ( \233 , \172 , \169 );
nand \g11981/U$1 ( \234 , \232 , \233 );
not \mul_6_19_g11492/U$4 ( \235 , \234 );
and \mul_6_19_g11492/U$2 ( \236 , \230 , \235 );
not \mul_6_19_g11528/U$1 ( \237 , \228 );
and \mul_6_19_g11492/U$5 ( \238 , \234 , \237 );
nor \mul_6_19_g11492/U$1 ( \239 , \236 , \238 );
not \mul_6_19_g11467/U$3 ( \240 , \239 );
nand \mul_6_19_g11720/U$1 ( \241 , \153 , \B[5] );
nand \mul_6_19_g11686/U$1 ( \242 , \79 , \B[4] );
xor \mul_6_19_g11516/U$1 ( \243 , \241 , \242 );
nand \mul_6_19_g11625/U$1 ( \244 , \136 , \B[7] );
xor \mul_6_19_g11516/U$1_r1 ( \245 , \243 , \244 );
not \mul_6_19_g11514/U$1 ( \246 , \245 );
not \mul_6_19_g11467/U$4 ( \247 , \246 );
or \mul_6_19_g11467/U$2 ( \248 , \240 , \247 );
not \mul_6_19_g11775/U$2 ( \249 , \239 );
nand \mul_6_19_g11775/U$1 ( \250 , \249 , \245 );
nand \mul_6_19_g11467/U$1 ( \251 , \248 , \250 );
xnor \mul_6_19_g11402/U$1_r1 ( \252 , \220 , \251 );
not \mul_6_19_g11340/U$4 ( \253 , \252 );
or \mul_6_19_g11340/U$2 ( \254 , \194 , \253 );
xor \mul_6_19_g11439/U$1 ( \255 , \201 , \208 );
xor \mul_6_19_g11439/U$1_r1 ( \256 , \255 , \216 );
xor \mul_6_19_g11510/U$1 ( \257 , \202 , \203 );
xor \mul_6_19_g11510/U$1_r1 ( \258 , \257 , \205 );
not \g11949/U$2 ( \259 , \258 );
nand \mul_6_19_g11717/U$1 ( \260 , \136 , \B[4] );
not \mul_6_19_g11560/U$3 ( \261 , \260 );
nand \mul_6_19_g11934/U$1 ( \262 , \104 , \B[8] );
not \mul_6_19_g11560/U$4 ( \263 , \262 );
or \mul_6_19_g11560/U$2 ( \264 , \261 , \263 );
and \mul_6_19_g11693/U$1 ( \265 , \111 , \B[9] );
nand \mul_6_19_g11560/U$1 ( \266 , \264 , \265 );
not \mul_6_19_g11788/U$2 ( \267 , \260 );
not \mul_6_19_g11734/U$1 ( \268 , \262 );
nand \mul_6_19_g11788/U$1 ( \269 , \267 , \268 );
nand \mul_6_19_g11534/U$1 ( \270 , \266 , \269 );
nand \g11949/U$1 ( \271 , \259 , \270 );
not \mul_6_19_g11517/U$1 ( \272 , \270 );
not \mul_6_19_g11482/U$3 ( \273 , \272 );
not \mul_6_19_g11482/U$4 ( \274 , \258 );
or \mul_6_19_g11482/U$2 ( \275 , \273 , \274 );
nand \mul_6_19_g11650/U$1 ( \276 , \95 , \B[5] );
not \mul_6_19_g11562/U$3 ( \277 , \276 );
nand \mul_6_19_g11632/U$1 ( \278 , \86 , \B[3] );
not \mul_6_19_g11562/U$4 ( \279 , \278 );
or \mul_6_19_g11562/U$2 ( \280 , \277 , \279 );
nand \mul_6_19_g11867/U$1 ( \281 , \127 , \B[6] );
not \mul_6_19_g11640/U$1 ( \282 , \281 );
nand \mul_6_19_g11562/U$1 ( \283 , \280 , \282 );
or \mul_6_19_g11781/U$1 ( \284 , \278 , \276 );
nand \mul_6_19_g11535/U$1 ( \285 , \283 , \284 );
nand \mul_6_19_g11482/U$1 ( \286 , \275 , \285 );
and \g11936/U$1 ( \287 , \271 , \286 );
xor \mul_6_19_g11394/U$4 ( \288 , \256 , \287 );
xor \mul_6_19_g11532/U$1 ( \289 , \210 , \211 );
xor \mul_6_19_g11532/U$1_r1 ( \290 , \289 , \213 );
xor \mul_6_19_g11519/U$1 ( \291 , \180 , \181 );
xor \mul_6_19_g11519/U$1_r1 ( \292 , \291 , \185 );
xor \mul_6_19_g11430/U$4 ( \293 , \290 , \292 );
nand \mul_6_19_g11694/U$1 ( \294 , \200 , \B[7] );
nand \mul_6_19_g11721/U$1 ( \295 , \79 , \B[0] );
not \mul_6_19_g11606/U$2 ( \296 , \295 );
and \mul_6_19_g11695/U$1 ( \297 , \152 , \B[1] );
nand \mul_6_19_g11606/U$1 ( \298 , \296 , \297 );
xor \mul_6_19_g11487/U$4 ( \299 , \294 , \298 );
xnor \g11818/U$1 ( \300 , \184 , \183 );
and \mul_6_19_g11487/U$3 ( \301 , \299 , \300 );
and \mul_6_19_g11487/U$5 ( \302 , \294 , \298 );
or \mul_6_19_g11487/U$2 ( \303 , \301 , \302 );
and \mul_6_19_g11430/U$3 ( \304 , \293 , \303 );
and \mul_6_19_g11430/U$5 ( \305 , \290 , \292 );
or \mul_6_19_g11430/U$2 ( \306 , \304 , \305 );
and \mul_6_19_g11394/U$3 ( \307 , \288 , \306 );
and \mul_6_19_g11394/U$5 ( \308 , \256 , \287 );
or \mul_6_19_g11394/U$2 ( \309 , \307 , \308 );
not \mul_6_19_g11393/U$1 ( \310 , \309 );
nand \mul_6_19_g11340/U$1 ( \311 , \254 , \310 );
or \g11944/U$1 ( \312 , \252 , \193 );
nand \mul_6_19_g11332/U$1 ( \313 , \311 , \312 );
nand \mul_6_19_g11497/U$1 ( \314 , \245 , \237 );
not \mul_6_19_g2/U$3 ( \315 , \314 );
not \mul_6_19_g2/U$4 ( \316 , \234 );
or \mul_6_19_g2/U$2 ( \317 , \315 , \316 );
or \mul_6_19_g2/U$5 ( \318 , \245 , \237 );
nand \mul_6_19_g2/U$1 ( \319 , \317 , \318 );
nand \mul_6_19_g11672/U$1 ( \320 , \136 , \B[8] );
nand \mul_6_19_g11636/U$1 ( \321 , \79 , \B[5] );
xor \mul_6_19_g11513/U$1 ( \322 , \320 , \321 );
nand \mul_6_19_g11685/U$1 ( \323 , \153 , \B[6] );
xor \mul_6_19_g11513/U$1_r1 ( \324 , \322 , \323 );
xor \mul_6_19_g11516/U$4 ( \325 , \241 , \242 );
and \mul_6_19_g11516/U$3 ( \326 , \325 , \244 );
and \mul_6_19_g11516/U$5 ( \327 , \241 , \242 );
or \mul_6_19_g11516/U$2 ( \328 , \326 , \327 );
and \mul_6_19_g11493/U$2 ( \329 , \324 , \328 );
not \mul_6_19_g11493/U$4 ( \330 , \324 );
not \mul_6_19_g11515/U$1 ( \331 , \328 );
and \mul_6_19_g11493/U$3 ( \332 , \330 , \331 );
nor \mul_6_19_g11493/U$1 ( \333 , \329 , \332 );
nand \mul_6_19_g11737/U$1 ( \334 , \95 , \B[9] );
nand \mul_6_19_g11747/U$1 ( \335 , \86 , \B[7] );
xor \mul_6_19_g11474/U$1 ( \336 , \334 , \335 );
xor \mul_6_19_g11512/U$4 ( \337 , \195 , \196 );
and \mul_6_19_g11512/U$3 ( \338 , \337 , \198 );
and \mul_6_19_g11512/U$5 ( \339 , \195 , \196 );
or \mul_6_19_g11512/U$2 ( \340 , \338 , \339 );
xor \mul_6_19_g11474/U$1_r1 ( \341 , \336 , \340 );
and \mul_6_19_g11449/U$2 ( \342 , \333 , \341 );
not \mul_6_19_g11449/U$4 ( \343 , \333 );
not \fopt11848/U$1 ( \344 , \341 );
and \mul_6_19_g11449/U$3 ( \345 , \343 , \344 );
or \mul_6_19_g11449/U$1 ( \346 , \342 , \345 );
xor \mul_6_19_g11355/U$1 ( \347 , \319 , \346 );
not \mul_6_19_g11415/U$3 ( \348 , \199 );
not \mul_6_19_g11442/U$1 ( \349 , \251 );
not \mul_6_19_g11415/U$4 ( \350 , \349 );
or \mul_6_19_g11415/U$2 ( \351 , \348 , \350 );
not \mul_6_19_g11438/U$1 ( \352 , \219 );
nand \mul_6_19_g11415/U$1 ( \353 , \351 , \352 );
not \mul_6_19_g11420/U$2 ( \354 , \199 );
nand \mul_6_19_g11420/U$1 ( \355 , \354 , \251 );
nand \mul_6_19_g11404/U$1 ( \356 , \353 , \355 );
xor \mul_6_19_g11355/U$1_r1 ( \357 , \347 , \356 );
or \mul_6_19_g11764/U$1 ( \358 , \313 , \357 );
xor \mul_6_19_g11474/U$4 ( \359 , \334 , \335 );
and \mul_6_19_g11474/U$3 ( \360 , \359 , \340 );
and \mul_6_19_g11474/U$5 ( \361 , \334 , \335 );
or \mul_6_19_g11474/U$2 ( \362 , \360 , \361 );
nand \mul_6_19_g11633/U$1 ( \363 , \86 , \B[8] );
xor \mul_6_19_g11513/U$4 ( \364 , \320 , \321 );
and \mul_6_19_g11513/U$3 ( \365 , \364 , \323 );
and \mul_6_19_g11513/U$5 ( \366 , \320 , \321 );
or \mul_6_19_g11513/U$2 ( \367 , \365 , \366 );
xor \mul_6_19_g11440/U$1 ( \368 , \363 , \367 );
nand \mul_6_19_g11749/U$1 ( \369 , \153 , \B[7] );
nand \mul_6_19_g11637/U$1 ( \370 , \79 , \B[6] );
xor \mul_6_19_g11530/U$1 ( \371 , \369 , \370 );
nand \mul_6_19_g11719/U$1 ( \372 , \136 , \B[9] );
xor \mul_6_19_g11530/U$1_r1 ( \373 , \371 , \372 );
xor \mul_6_19_g11440/U$1_r1 ( \374 , \368 , \373 );
xor \mul_6_19_g11371/U$1 ( \375 , \362 , \374 );
nand \mul_6_19_g11450/U$1 ( \376 , \341 , \324 );
and \mul_6_19_g11425/U$2 ( \377 , \376 , \331 );
nor \mul_6_19_g11455/U$1 ( \378 , \341 , \324 );
nor \mul_6_19_g11425/U$1 ( \379 , \377 , \378 );
xor \mul_6_19_g11371/U$1_r1 ( \380 , \375 , \379 );
not \mul_6_19_g11768/U$2 ( \381 , \380 );
xor \mul_6_19_g11355/U$4 ( \382 , \319 , \346 );
and \mul_6_19_g11355/U$3 ( \383 , \382 , \356 );
and \mul_6_19_g11355/U$5 ( \384 , \319 , \346 );
or \mul_6_19_g11355/U$2 ( \385 , \383 , \384 );
nor \mul_6_19_g11768/U$1 ( \386 , \381 , \385 );
not \fopt11898/U$1 ( \387 , \386 );
nand \mul_6_19_g11858/U$1 ( \388 , \358 , \387 );
xor \mul_6_19_g11530/U$4 ( \389 , \369 , \370 );
and \mul_6_19_g11530/U$3 ( \390 , \389 , \372 );
and \mul_6_19_g11530/U$5 ( \391 , \369 , \370 );
or \mul_6_19_g11530/U$2 ( \392 , \390 , \391 );
xor \mul_6_19_g11520/U$1 ( \393 , \156 , \157 );
xor \mul_6_19_g11520/U$1_r1 ( \394 , \393 , \159 );
xor \mul_6_19_g11407/U$4 ( \395 , \392 , \394 );
xor \mul_6_19_g11440/U$4 ( \396 , \363 , \367 );
and \mul_6_19_g11440/U$3 ( \397 , \396 , \373 );
and \mul_6_19_g11440/U$5 ( \398 , \363 , \367 );
or \mul_6_19_g11440/U$2 ( \399 , \397 , \398 );
and \mul_6_19_g11407/U$3 ( \400 , \395 , \399 );
and \mul_6_19_g11407/U$5 ( \401 , \392 , \394 );
or \mul_6_19_g11407/U$2 ( \402 , \400 , \401 );
xor \mul_6_19_g11476/U$1 ( \403 , \147 , \154 );
xor \mul_6_19_g11476/U$1_r1 ( \404 , \403 , \162 );
nand \mul_6_19_g11395/U$1 ( \405 , \402 , \404 );
xor \mul_6_19_g11371/U$4 ( \406 , \362 , \374 );
and \mul_6_19_g11371/U$3 ( \407 , \406 , \379 );
and \mul_6_19_g11371/U$5 ( \408 , \362 , \374 );
or \mul_6_19_g11371/U$2 ( \409 , \407 , \408 );
xor \mul_6_19_g11407/U$1 ( \410 , \392 , \394 );
xor \mul_6_19_g11407/U$1_r1 ( \411 , \410 , \399 );
nand \mul_6_19_g11357/U$1 ( \412 , \409 , \411 );
nand \mul_6_19_g11344/U$1 ( \413 , \405 , \412 );
nor \mul_6_19_g11277/U$1 ( \414 , \388 , \413 );
not \mul_6_19_g11762/U$2 ( \415 , \414 );
xor \mul_6_19_g11394/U$1 ( \416 , \256 , \287 );
xor \mul_6_19_g11394/U$1_r1 ( \417 , \416 , \306 );
xor \mul_6_19_g11475/U$1 ( \418 , \190 , \191 );
and \mul_6_19_g11436/U$2 ( \419 , \418 , \188 );
not \mul_6_19_g11436/U$4 ( \420 , \418 );
not \mul_6_19_g11518/U$1 ( \421 , \188 );
and \mul_6_19_g11436/U$3 ( \422 , \420 , \421 );
or \mul_6_19_g11436/U$1 ( \423 , \419 , \422 );
xor \g11855/U$1 ( \424 , \417 , \423 );
not \mul_6_19_g11494/U$3 ( \425 , \285 );
not \mul_6_19_g11494/U$4 ( \426 , \272 );
or \mul_6_19_g11494/U$2 ( \427 , \425 , \426 );
not \mul_6_19_g11776/U$2 ( \428 , \285 );
nand \mul_6_19_g11776/U$1 ( \429 , \428 , \270 );
nand \mul_6_19_g11494/U$1 ( \430 , \427 , \429 );
and \mul_6_19_g11466/U$2 ( \431 , \430 , \258 );
not \mul_6_19_g11466/U$4 ( \432 , \430 );
not \fopt11895/U$1 ( \433 , \258 );
and \mul_6_19_g11466/U$3 ( \434 , \432 , \433 );
nor \mul_6_19_g11466/U$1 ( \435 , \431 , \434 );
nand \mul_6_19_g11758/U$1 ( \436 , \95 , \B[4] );
nand \mul_6_19_g11663/U$1 ( \437 , \86 , \B[2] );
xor \mul_6_19_g11556/U$4 ( \438 , \436 , \437 );
nand \mul_6_19_g11664/U$1 ( \439 , \B[9] , \118 );
and \mul_6_19_g11556/U$3 ( \440 , \438 , \439 );
and \mul_6_19_g11556/U$5 ( \441 , \436 , \437 );
or \mul_6_19_g11556/U$2 ( \442 , \440 , \441 );
xor \mul_6_19_g11759/U$1 ( \443 , \276 , \281 );
xor \mul_6_19_g11759/U$1_r1 ( \444 , \443 , \278 );
xor \mul_6_19_g11445/U$4 ( \445 , \442 , \444 );
and \mul_6_19_g11711/U$1 ( \446 , \136 , \B[3] );
and \mul_6_19_g11708/U$1 ( \447 , \104 , \B[7] );
or \mul_6_19_g11787/U$1 ( \448 , \446 , \447 );
nand \mul_6_19_g11671/U$1 ( \449 , \111 , \B[8] );
not \mul_6_19_g11670/U$1 ( \450 , \449 );
and \mul_6_19_g11537/U$2 ( \451 , \448 , \450 );
and \mul_6_19_g11576/U$2 ( \452 , \446 , \447 );
nor \mul_6_19_g11537/U$1 ( \453 , \451 , \452 );
and \mul_6_19_g11445/U$3 ( \454 , \445 , \453 );
and \mul_6_19_g11445/U$5 ( \455 , \442 , \444 );
or \mul_6_19_g11445/U$2 ( \456 , \454 , \455 );
xor \mul_6_19_g11373/U$4 ( \457 , \435 , \456 );
xor \g11811/U$1 ( \458 , \260 , \268 );
xor \g11811/U$1_r1 ( \459 , \458 , \265 );
nand \mul_6_19_g11626/U$1 ( \460 , \200 , \B[6] );
nand \mul_6_19_g11643/U$1 ( \461 , \127 , \B[5] );
xor \mul_6_19_g11507/U$4 ( \462 , \460 , \461 );
not \mul_6_19_g11593/U$3 ( \463 , \297 );
not \mul_6_19_g11593/U$4 ( \464 , \295 );
and \mul_6_19_g11593/U$2 ( \465 , \463 , \464 );
and \mul_6_19_g11593/U$5 ( \466 , \297 , \295 );
nor \mul_6_19_g11593/U$1 ( \467 , \465 , \466 );
and \mul_6_19_g11507/U$3 ( \468 , \462 , \467 );
and \mul_6_19_g11507/U$5 ( \469 , \460 , \461 );
or \mul_6_19_g11507/U$2 ( \470 , \468 , \469 );
xor \mul_6_19_g11418/U$4 ( \471 , \459 , \470 );
and \mul_6_19_g11677/U$1 ( \472 , \86 , \B[0] );
nand \mul_6_19_g11612/U$1 ( \473 , \297 , \472 );
nand \mul_6_19_g11683/U$1 ( \474 , \143 , \B[5] );
not \mul_6_19_g11582/U$3 ( \475 , \474 );
nand \mul_6_19_g11700/U$1 ( \476 , \127 , \B[4] );
not \mul_6_19_g11582/U$4 ( \477 , \476 );
or \mul_6_19_g11582/U$2 ( \478 , \475 , \477 );
and \mul_6_19_g11738/U$1 ( \479 , \136 , \B[2] );
nand \mul_6_19_g11582/U$1 ( \480 , \478 , \479 );
not \mul_6_19_g11599/U$2 ( \481 , \476 );
not \mul_6_19_g11682/U$1 ( \482 , \474 );
nand \mul_6_19_g11599/U$1 ( \483 , \481 , \482 );
nand \mul_6_19_g11571/U$1 ( \484 , \480 , \483 );
not \mul_6_19_g11549/U$1 ( \485 , \484 );
xor \mul_6_19_g11463/U$4 ( \486 , \473 , \485 );
nand \mul_6_19_g11752/U$1 ( \487 , \111 , \B[7] );
nand \mul_6_19_g11673/U$1 ( \488 , \95 , \B[3] );
nand \mul_6_19_g11616/U$1 ( \489 , \487 , \488 );
and \mul_6_19_g11648/U$1 ( \490 , \118 , \B[8] );
and \mul_6_19_g11538/U$2 ( \491 , \489 , \490 );
nor \mul_6_19_g11614/U$1 ( \492 , \487 , \488 );
nor \mul_6_19_g11538/U$1 ( \493 , \491 , \492 );
and \mul_6_19_g11463/U$3 ( \494 , \486 , \493 );
and \mul_6_19_g11463/U$5 ( \495 , \473 , \485 );
or \mul_6_19_g11463/U$2 ( \496 , \494 , \495 );
and \mul_6_19_g11418/U$3 ( \497 , \471 , \496 );
and \mul_6_19_g11418/U$5 ( \498 , \459 , \470 );
or \mul_6_19_g11418/U$2 ( \499 , \497 , \498 );
and \mul_6_19_g11373/U$3 ( \500 , \457 , \499 );
and \mul_6_19_g11373/U$5 ( \501 , \435 , \456 );
or \mul_6_19_g11373/U$2 ( \502 , \500 , \501 );
xnor \mul_6_19_g11334/U$1 ( \503 , \424 , \502 );
xor \mul_6_19_g11430/U$1 ( \504 , \290 , \292 );
xor \mul_6_19_g11430/U$1_r1 ( \505 , \504 , \303 );
xor \mul_6_19_g11487/U$1 ( \506 , \294 , \298 );
xor \mul_6_19_g11487/U$1_r1 ( \507 , \506 , \300 );
xor \mul_6_19_g11445/U$1 ( \508 , \442 , \444 );
xor \mul_6_19_g11445/U$1_r1 ( \509 , \508 , \453 );
xor \mul_6_19_g11375/U$4 ( \510 , \507 , \509 );
xor \mul_6_19_g11576/U$1 ( \511 , \446 , \447 );
and \mul_6_19_g11547/U$2 ( \512 , \511 , \450 );
not \mul_6_19_g11547/U$4 ( \513 , \511 );
and \mul_6_19_g11547/U$3 ( \514 , \513 , \449 );
nor \mul_6_19_g11547/U$1 ( \515 , \512 , \514 );
not \mul_6_19_g11531/U$1 ( \516 , \515 );
xor \mul_6_19_g11556/U$1 ( \517 , \436 , \437 );
xor \mul_6_19_g11556/U$1_r1 ( \518 , \517 , \439 );
nand \mul_6_19_g11502/U$1 ( \519 , \516 , \518 );
and \mul_6_19_g11696/U$1 ( \520 , \104 , \B[6] );
and \mul_6_19_g11638/U$1 ( \521 , \86 , \B[1] );
not \mul_6_19_g11594/U$3 ( \522 , \521 );
nand \mul_6_19_g11733/U$1 ( \523 , \153 , \B[0] );
not \mul_6_19_g11594/U$4 ( \524 , \523 );
or \mul_6_19_g11594/U$2 ( \525 , \522 , \524 );
or \mul_6_19_g11594/U$5 ( \526 , \521 , \523 );
nand \mul_6_19_g11594/U$1 ( \527 , \525 , \526 );
xor \mul_6_19_g11486/U$4 ( \528 , \520 , \527 );
and \mul_6_19_g11741/U$1 ( \529 , \136 , \B[1] );
and \mul_6_19_g11575/U$2 ( \530 , \472 , \529 );
and \mul_6_19_g11486/U$3 ( \531 , \528 , \530 );
and \mul_6_19_g11486/U$5 ( \532 , \520 , \527 );
or \mul_6_19_g11486/U$2 ( \533 , \531 , \532 );
and \mul_6_19_g11434/U$2 ( \534 , \519 , \533 );
nor \mul_6_19_g11501/U$1 ( \535 , \516 , \518 );
nor \mul_6_19_g11434/U$1 ( \536 , \534 , \535 );
and \mul_6_19_g11375/U$3 ( \537 , \510 , \536 );
and \mul_6_19_g11375/U$5 ( \538 , \507 , \509 );
or \mul_6_19_g11375/U$2 ( \539 , \537 , \538 );
xor \mul_6_19_g11879/U$4 ( \540 , \505 , \539 );
xor \mul_6_19_g11373/U$1 ( \541 , \435 , \456 );
xor \mul_6_19_g11373/U$1_r1 ( \542 , \541 , \499 );
and \mul_6_19_g11879/U$3 ( \543 , \540 , \542 );
and \mul_6_19_g11879/U$5 ( \544 , \505 , \539 );
or \mul_6_19_g11879/U$2 ( \545 , \543 , \544 );
nand \mul_6_19_g11309/U$1 ( \546 , \503 , \545 );
not \mul_6_19_g11339/U$3 ( \547 , \417 );
not \mul_6_19_g11427/U$1 ( \548 , \423 );
not \mul_6_19_g11339/U$4 ( \549 , \548 );
or \mul_6_19_g11339/U$2 ( \550 , \547 , \549 );
not \mul_6_19_g11372/U$1 ( \551 , \502 );
nand \mul_6_19_g11339/U$1 ( \552 , \550 , \551 );
not \mul_6_19_g11769/U$2 ( \553 , \417 );
nand \mul_6_19_g11769/U$1 ( \554 , \553 , \423 );
nand \mul_6_19_g11331/U$1 ( \555 , \552 , \554 );
not \mul_6_19_g11765/U$2 ( \556 , \555 );
xor \mul_6_19_g11841/U$1 ( \557 , \193 , \309 );
xor \mul_6_19_g11841/U$1_r1 ( \558 , \557 , \252 );
nand \mul_6_19_g11765/U$1 ( \559 , \556 , \558 );
nand \mul_6_19_g11294/U$1 ( \560 , \546 , \559 );
nor \mul_6_19_g11762/U$1 ( \561 , \415 , \560 );
not \mul_6_19_g11249/U$3 ( \562 , \561 );
nand \mul_6_19_g11657/U$1 ( \563 , \136 , \B[0] );
not \mul_6_19_g11590/U$3 ( \564 , \563 );
and \mul_6_19_g11623/U$1 ( \565 , \95 , \B[1] );
not \mul_6_19_g11590/U$4 ( \566 , \565 );
and \mul_6_19_g11590/U$2 ( \567 , \564 , \566 );
and \mul_6_19_g11590/U$5 ( \568 , \563 , \565 );
nor \mul_6_19_g11590/U$1 ( \569 , \567 , \568 );
nand \mul_6_19_g11736/U$1 ( \570 , \111 , \B[4] );
nand \mul_6_19_g11624/U$1 ( \571 , \200 , \B[2] );
xor \mul_6_19_g11550/U$4 ( \572 , \570 , \571 );
nand \mul_6_19_g11743/U$1 ( \573 , \104 , \B[3] );
and \mul_6_19_g11550/U$3 ( \574 , \572 , \573 );
and \mul_6_19_g11550/U$5 ( \575 , \570 , \571 );
or \mul_6_19_g11550/U$2 ( \576 , \574 , \575 );
xor \mul_6_19_g11465/U$4 ( \577 , \569 , \576 );
nand \mul_6_19_g11654/U$1 ( \578 , \104 , \B[4] );
and \mul_6_19_g11760/U$1 ( \579 , \143 , \B[3] );
xor \g12010/U$1 ( \580 , \578 , \579 );
nand \mul_6_19_g11732/U$1 ( \581 , \127 , \B[2] );
xnor \g12010/U$1_r1 ( \582 , \580 , \581 );
and \mul_6_19_g11465/U$3 ( \583 , \577 , \582 );
and \mul_6_19_g11465/U$5 ( \584 , \569 , \576 );
or \mul_6_19_g11465/U$2 ( \585 , \583 , \584 );
not \mul_6_19_g11426/U$3 ( \586 , \585 );
not \mul_6_19_g11780/U$2 ( \587 , \565 );
nor \mul_6_19_g11780/U$1 ( \588 , \587 , \563 );
xor \mul_6_19_g11575/U$1 ( \589 , \472 , \529 );
xor \mul_6_19_g11478/U$1 ( \590 , \588 , \589 );
not \mul_6_19_g11583/U$3 ( \591 , \581 );
not \mul_6_19_g11583/U$4 ( \592 , \578 );
or \mul_6_19_g11583/U$2 ( \593 , \591 , \592 );
nand \mul_6_19_g11583/U$1 ( \594 , \593 , \579 );
or \mul_6_19_g11783/U$1 ( \595 , \578 , \581 );
nand \mul_6_19_g11572/U$1 ( \596 , \594 , \595 );
xor \mul_6_19_g11478/U$1_r1 ( \597 , \590 , \596 );
not \mul_6_19_g11426/U$4 ( \598 , \597 );
and \mul_6_19_g11426/U$2 ( \599 , \586 , \598 );
and \mul_6_19_g11426/U$5 ( \600 , \585 , \597 );
nor \mul_6_19_g11426/U$1 ( \601 , \599 , \600 );
nand \mul_6_19_g11628/U$1 ( \602 , \95 , \B[2] );
nand \mul_6_19_g11740/U$1 ( \603 , \104 , \B[5] );
xor \mul_6_19_g11789/U$1 ( \604 , \602 , \603 );
nand \mul_6_19_g11666/U$1 ( \605 , \111 , \B[6] );
xor \mul_6_19_g11789/U$1_r1 ( \606 , \604 , \605 );
not \mul_6_19_g11553/U$1 ( \607 , \606 );
not \mul_6_19_g11503/U$3 ( \608 , \607 );
nand \mul_6_19_g11669/U$1 ( \609 , \118 , \B[7] );
and \g11988/U$1 ( \610 , \127 , \B[3] );
xor \g11957/U$1 ( \611 , \609 , \610 );
nand \mul_6_19_g11748/U$1 ( \612 , \200 , \B[4] );
xnor \g11957/U$1_r1 ( \613 , \611 , \612 );
not \mul_6_19_g11503/U$4 ( \614 , \613 );
or \mul_6_19_g11503/U$2 ( \615 , \608 , \614 );
not \mul_6_19_g11551/U$1 ( \616 , \613 );
nand \mul_6_19_g11504/U$1 ( \617 , \616 , \606 );
nand \mul_6_19_g11503/U$1 ( \618 , \615 , \617 );
and \mul_6_19_g11725/U$1 ( \619 , \118 , \B[6] );
not \mul_6_19_g11724/U$1 ( \620 , \619 );
nand \mul_6_19_g11704/U$1 ( \621 , \111 , \B[5] );
or \mul_6_19_g11540/U$2 ( \622 , \620 , \621 );
not \mul_6_19_g11563/U$3 ( \623 , \621 );
not \mul_6_19_g11563/U$4 ( \624 , \620 );
or \mul_6_19_g11563/U$2 ( \625 , \623 , \624 );
nand \mul_6_19_g11661/U$1 ( \626 , \127 , \B[1] );
not \mul_6_19_g11608/U$2 ( \627 , \626 );
and \mul_6_19_g11713/U$1 ( \628 , \95 , \B[0] );
nand \mul_6_19_g11608/U$1 ( \629 , \627 , \628 );
not \mul_6_19_g11577/U$1 ( \630 , \629 );
nand \mul_6_19_g11563/U$1 ( \631 , \625 , \630 );
nand \mul_6_19_g11540/U$1 ( \632 , \622 , \631 );
not \mul_6_19_g11511/U$1 ( \633 , \632 );
and \mul_6_19_g11461/U$2 ( \634 , \618 , \633 );
not \mul_6_19_g11461/U$4 ( \635 , \618 );
and \mul_6_19_g11461/U$3 ( \636 , \635 , \632 );
nor \mul_6_19_g11461/U$1 ( \637 , \634 , \636 );
not \mul_6_19_g11444/U$1 ( \638 , \637 );
and \mul_6_19_g11405/U$2 ( \639 , \601 , \638 );
not \mul_6_19_g11405/U$4 ( \640 , \601 );
and \mul_6_19_g11405/U$3 ( \641 , \640 , \637 );
nor \mul_6_19_g11405/U$1 ( \642 , \639 , \641 );
xor \g11815/U$1 ( \643 , \619 , \621 );
xnor \g11815/U$1_r1 ( \644 , \643 , \629 );
nand \mul_6_19_g11726/U$1 ( \645 , \118 , \B[5] );
nand \mul_6_19_g11698/U$1 ( \646 , \127 , \B[0] );
not \mul_6_19_g11613/U$2 ( \647 , \646 );
and \mul_6_19_g11761/U$1 ( \648 , \143 , \B[1] );
nand \mul_6_19_g11613/U$1 ( \649 , \647 , \648 );
xor \mul_6_19_g11489/U$4 ( \650 , \645 , \649 );
not \mul_6_19_g11588/U$3 ( \651 , \628 );
not \mul_6_19_g11588/U$4 ( \652 , \626 );
and \mul_6_19_g11588/U$2 ( \653 , \651 , \652 );
and \mul_6_19_g11588/U$5 ( \654 , \626 , \628 );
nor \mul_6_19_g11588/U$1 ( \655 , \653 , \654 );
and \mul_6_19_g11489/U$3 ( \656 , \650 , \655 );
and \mul_6_19_g11489/U$5 ( \657 , \645 , \649 );
or \mul_6_19_g11489/U$2 ( \658 , \656 , \657 );
xor \mul_6_19_g11412/U$4 ( \659 , \644 , \658 );
xor \mul_6_19_g11465/U$1 ( \660 , \569 , \576 );
xor \mul_6_19_g11465/U$1_r1 ( \661 , \660 , \582 );
and \mul_6_19_g11412/U$3 ( \662 , \659 , \661 );
and \mul_6_19_g11412/U$5 ( \663 , \644 , \658 );
or \mul_6_19_g11412/U$2 ( \664 , \662 , \663 );
nand \mul_6_19_g11381/U$1 ( \665 , \642 , \664 );
not \mul_6_19_g11320/U$3 ( \666 , \665 );
xor \mul_6_19_g11412/U$1 ( \667 , \644 , \658 );
xor \mul_6_19_g11412/U$1_r1 ( \668 , \667 , \661 );
nand \mul_6_19_g11642/U$1 ( \669 , \118 , \B[4] );
nand \mul_6_19_g11678/U$1 ( \670 , \104 , \B[2] );
xor \mul_6_19_g11557/U$4 ( \671 , \669 , \670 );
nand \mul_6_19_g11639/U$1 ( \672 , \111 , \B[3] );
and \mul_6_19_g11557/U$3 ( \673 , \671 , \672 );
and \mul_6_19_g11557/U$5 ( \674 , \669 , \670 );
or \mul_6_19_g11557/U$2 ( \675 , \673 , \674 );
xor \mul_6_19_g11550/U$1 ( \676 , \570 , \571 );
xor \mul_6_19_g11550/U$1_r1 ( \677 , \676 , \573 );
xor \mul_6_19_g11448/U$4 ( \678 , \675 , \677 );
xor \mul_6_19_g11489/U$1 ( \679 , \645 , \649 );
xor \mul_6_19_g11489/U$1_r1 ( \680 , \679 , \655 );
and \mul_6_19_g11448/U$3 ( \681 , \678 , \680 );
and \mul_6_19_g11448/U$5 ( \682 , \675 , \677 );
or \mul_6_19_g11448/U$2 ( \683 , \681 , \682 );
nand \mul_6_19_g11397/U$1 ( \684 , \668 , \683 );
not \mul_6_19_g11350/U$3 ( \685 , \684 );
xor \mul_6_19_g11448/U$1 ( \686 , \675 , \677 );
xor \mul_6_19_g11448/U$1_r1 ( \687 , \686 , \680 );
nand \mul_6_19_g11652/U$1 ( \688 , \200 , \B[0] );
not \mul_6_19_g11782/U$2 ( \689 , \688 );
and \mul_6_19_g11684/U$1 ( \690 , \104 , \B[1] );
nand \mul_6_19_g11782/U$1 ( \691 , \689 , \690 );
not \mul_6_19_g11591/U$3 ( \692 , \648 );
not \mul_6_19_g11591/U$4 ( \693 , \646 );
and \mul_6_19_g11591/U$2 ( \694 , \692 , \693 );
and \mul_6_19_g11591/U$5 ( \695 , \648 , \646 );
nor \mul_6_19_g11591/U$1 ( \696 , \694 , \695 );
xor \mul_6_19_g11481/U$4 ( \697 , \691 , \696 );
xor \mul_6_19_g11557/U$1 ( \698 , \669 , \670 );
xor \mul_6_19_g11557/U$1_r1 ( \699 , \698 , \672 );
and \mul_6_19_g11481/U$3 ( \700 , \697 , \699 );
and \mul_6_19_g11481/U$5 ( \701 , \691 , \696 );
or \mul_6_19_g11481/U$2 ( \702 , \700 , \701 );
nand \mul_6_19_g11423/U$1 ( \703 , \687 , \702 );
not \mul_6_19_g11385/U$3 ( \704 , \703 );
xor \mul_6_19_g11481/U$1 ( \705 , \691 , \696 );
xor \mul_6_19_g11481/U$1_r1 ( \706 , \705 , \699 );
not \mul_6_19_g11592/U$3 ( \707 , \690 );
not \mul_6_19_g11592/U$4 ( \708 , \688 );
and \mul_6_19_g11592/U$2 ( \709 , \707 , \708 );
and \mul_6_19_g11592/U$5 ( \710 , \688 , \690 );
nor \mul_6_19_g11592/U$1 ( \711 , \709 , \710 );
not \g11865/U$2 ( \712 , \711 );
and \mul_6_19_g11620/U$1 ( \713 , \118 , \B[3] );
not \g11866/U$2 ( \714 , \713 );
nand \mul_6_19_g11705/U$1 ( \715 , \111 , \B[2] );
nand \g11866/U$1 ( \716 , \714 , \715 );
nand \g11865/U$1 ( \717 , \712 , \716 );
not \mul_6_19_g11607/U$2 ( \718 , \715 );
nand \mul_6_19_g11607/U$1 ( \719 , \718 , \713 );
and \mul_6_19_g11539/U$1 ( \720 , \717 , \719 );
or \mul_6_19_g11773/U$1 ( \721 , \706 , \720 );
and \mul_6_19_g11729/U$1 ( \722 , \104 , \B[0] );
and \mul_6_19_g11646/U$1 ( \723 , \118 , \B[2] );
and \mul_6_19_g11574/U$2 ( \724 , \722 , \723 );
not \mul_6_19_g11779/U$2 ( \725 , \724 );
not \mul_6_19_g11546/U$3 ( \726 , \711 );
not \mul_6_19_g11597/U$3 ( \727 , \715 );
not \mul_6_19_g11597/U$4 ( \728 , \713 );
or \mul_6_19_g11597/U$2 ( \729 , \727 , \728 );
or \mul_6_19_g11597/U$5 ( \730 , \713 , \715 );
nand \mul_6_19_g11597/U$1 ( \731 , \729 , \730 );
not \mul_6_19_g11546/U$4 ( \732 , \731 );
and \mul_6_19_g11546/U$2 ( \733 , \726 , \732 );
and \mul_6_19_g11546/U$5 ( \734 , \731 , \711 );
nor \mul_6_19_g11546/U$1 ( \735 , \733 , \734 );
nand \mul_6_19_g11779/U$1 ( \736 , \725 , \735 );
not \g11955/U$3 ( \737 , \736 );
nand \mul_6_19_g11691/U$1 ( \738 , \111 , \B[1] );
not \mul_6_19_g11690/U$1 ( \739 , \738 );
nand \mul_6_19_g11645/U$1 ( \740 , \118 , \B[0] );
nor \mul_6_19_g11615/U$1 ( \741 , \738 , \740 );
xor \mul_6_19_g11484/U$4 ( \742 , \739 , \741 );
xor \mul_6_19_g11574/U$1 ( \743 , \722 , \723 );
and \mul_6_19_g11484/U$3 ( \744 , \742 , \743 );
and \mul_6_19_g11484/U$5 ( \745 , \739 , \741 );
or \mul_6_19_g11484/U$2 ( \746 , \744 , \745 );
not \g11955/U$4 ( \747 , \746 );
or \g11955/U$2 ( \748 , \737 , \747 );
not \mul_6_19_g11777/U$2 ( \749 , \735 );
nand \mul_6_19_g11777/U$1 ( \750 , \749 , \724 );
nand \g11955/U$1 ( \751 , \748 , \750 );
nand \mul_6_19_g11453/U$1 ( \752 , \706 , \720 );
nand \mul_6_19_g11424/U$1 ( \753 , \751 , \752 );
nand \mul_6_19_g11416/U$1 ( \754 , \721 , \753 );
not \mul_6_19_g11385/U$4 ( \755 , \754 );
or \mul_6_19_g11385/U$2 ( \756 , \704 , \755 );
or \mul_6_19_g11772/U$1 ( \757 , \687 , \702 );
nand \mul_6_19_g11385/U$1 ( \758 , \756 , \757 );
not \mul_6_19_g11350/U$4 ( \759 , \758 );
or \mul_6_19_g11350/U$2 ( \760 , \685 , \759 );
not \mul_6_19_g11410/U$1 ( \761 , \668 );
not \mul_6_19_g11447/U$1 ( \762 , \683 );
nand \mul_6_19_g11396/U$1 ( \763 , \761 , \762 );
nand \mul_6_19_g11350/U$1 ( \764 , \760 , \763 );
not \mul_6_19_g11320/U$4 ( \765 , \764 );
or \mul_6_19_g11320/U$2 ( \766 , \666 , \765 );
not \mul_6_19_g11400/U$1 ( \767 , \642 );
not \mul_6_19_g11411/U$1 ( \768 , \664 );
nand \mul_6_19_g11380/U$1 ( \769 , \767 , \768 );
nand \mul_6_19_g11320/U$1 ( \770 , \766 , \769 );
not \mul_6_19_g11470/U$3 ( \771 , \606 );
not \mul_6_19_g11470/U$4 ( \772 , \613 );
or \mul_6_19_g11470/U$2 ( \773 , \771 , \772 );
nand \mul_6_19_g11470/U$1 ( \774 , \773 , \632 );
nand \mul_6_19_g11505/U$1 ( \775 , \616 , \607 );
nand \mul_6_19_g11458/U$1 ( \776 , \774 , \775 );
not \mul_6_19_g11581/U$3 ( \777 , \612 );
not \mul_6_19_g11581/U$4 ( \778 , \609 );
or \mul_6_19_g11581/U$2 ( \779 , \777 , \778 );
nand \mul_6_19_g11581/U$1 ( \780 , \779 , \610 );
or \mul_6_19_g11786/U$1 ( \781 , \612 , \609 );
nand \mul_6_19_g11569/U$1 ( \782 , \780 , \781 );
not \mul_6_19_g11580/U$3 ( \783 , \603 );
not \mul_6_19_g11580/U$4 ( \784 , \605 );
or \mul_6_19_g11580/U$2 ( \785 , \783 , \784 );
not \mul_6_19_g11627/U$1 ( \786 , \602 );
nand \mul_6_19_g11580/U$1 ( \787 , \785 , \786 );
or \mul_6_19_g11785/U$1 ( \788 , \603 , \605 );
nand \mul_6_19_g11570/U$1 ( \789 , \787 , \788 );
xor \mul_6_19_g11488/U$1 ( \790 , \782 , \789 );
xor \g12023/U$1 ( \791 , \479 , \476 );
not \g12023/U$2 ( \792 , \474 );
xor \g12023/U$1_r1 ( \793 , \791 , \792 );
not \mul_6_19_g11548/U$1 ( \794 , \793 );
and \mul_6_19_g11462/U$2 ( \795 , \790 , \794 );
not \mul_6_19_g11462/U$4 ( \796 , \790 );
and \mul_6_19_g11462/U$3 ( \797 , \796 , \793 );
nor \mul_6_19_g11462/U$1 ( \798 , \795 , \797 );
xor \mul_6_19_g11379/U$1 ( \799 , \776 , \798 );
xor \mul_6_19_g11541/U$1 ( \800 , \488 , \487 );
xor \mul_6_19_g11541/U$1_r1 ( \801 , \800 , \490 );
xor \mul_6_19_g11486/U$1 ( \802 , \520 , \527 );
xor \mul_6_19_g11486/U$1_r1 ( \803 , \802 , \530 );
xor \mul_6_19_g11409/U$1 ( \804 , \801 , \803 );
xor \mul_6_19_g11478/U$4 ( \805 , \588 , \589 );
and \mul_6_19_g11478/U$3 ( \806 , \805 , \596 );
and \mul_6_19_g11478/U$5 ( \807 , \588 , \589 );
or \mul_6_19_g11478/U$2 ( \808 , \806 , \807 );
xor \mul_6_19_g11409/U$1_r1 ( \809 , \804 , \808 );
xor \mul_6_19_g11379/U$1_r1 ( \810 , \799 , \809 );
not \mul_6_19_g11377/U$1 ( \811 , \810 );
not \g11953/U$3 ( \812 , \597 );
not \g11953/U$4 ( \813 , \638 );
or \g11953/U$2 ( \814 , \812 , \813 );
not \mul_6_19_g11954/U$1 ( \815 , \597 );
not \mul_6_19_g11414/U$3 ( \816 , \815 );
not \mul_6_19_g11414/U$4 ( \817 , \637 );
or \mul_6_19_g11414/U$2 ( \818 , \816 , \817 );
not \mul_6_19_g11464/U$1 ( \819 , \585 );
nand \mul_6_19_g11414/U$1 ( \820 , \818 , \819 );
nand \g11953/U$1 ( \821 , \814 , \820 );
not \mul_6_19_g11401/U$1 ( \822 , \821 );
nand \mul_6_19_g11361/U$1 ( \823 , \811 , \822 );
nand \mul_6_19_g11285/U$1 ( \824 , \770 , \823 );
and \g12008/U$2 ( \825 , \518 , \515 );
not \g12008/U$4 ( \826 , \518 );
and \g12008/U$3 ( \827 , \826 , \516 );
or \g12008/U$1 ( \828 , \825 , \827 );
xor \mul_6_19_g11774/U$1 ( \829 , \828 , \533 );
xor \mul_6_19_g11409/U$4 ( \830 , \801 , \803 );
and \mul_6_19_g11409/U$3 ( \831 , \830 , \808 );
and \mul_6_19_g11409/U$5 ( \832 , \801 , \803 );
or \mul_6_19_g11409/U$2 ( \833 , \831 , \832 );
xor \mul_6_19_g11376/U$1 ( \834 , \829 , \833 );
xor \mul_6_19_g11507/U$1 ( \835 , \460 , \461 );
xor \mul_6_19_g11507/U$1_r1 ( \836 , \835 , \467 );
xor \mul_6_19_g11463/U$1 ( \837 , \473 , \485 );
xor \mul_6_19_g11463/U$1_r1 ( \838 , \837 , \493 );
xor \mul_6_19_g11391/U$1 ( \839 , \836 , \838 );
or \mul_6_19_g11778/U$1 ( \840 , \782 , \789 );
and \mul_6_19_g11457/U$2 ( \841 , \840 , \794 );
and \mul_6_19_g11488/U$2 ( \842 , \782 , \789 );
nor \mul_6_19_g11457/U$1 ( \843 , \841 , \842 );
xor \mul_6_19_g11391/U$1_r1 ( \844 , \839 , \843 );
not \mul_6_19_g11388/U$1 ( \845 , \844 );
and \mul_6_19_g11351/U$2 ( \846 , \834 , \845 );
not \mul_6_19_g11351/U$4 ( \847 , \834 );
and \mul_6_19_g11351/U$3 ( \848 , \847 , \844 );
nor \mul_6_19_g11351/U$1 ( \849 , \846 , \848 );
xor \mul_6_19_g11379/U$4 ( \850 , \776 , \798 );
and \mul_6_19_g11379/U$3 ( \851 , \850 , \809 );
and \mul_6_19_g11379/U$5 ( \852 , \776 , \798 );
or \mul_6_19_g11379/U$2 ( \853 , \851 , \852 );
nand \mul_6_19_g11327/U$1 ( \854 , \849 , \853 );
nand \mul_6_19_g11360/U$1 ( \855 , \810 , \821 );
and \mul_6_19_g11314/U$1 ( \856 , \854 , \855 );
nand \mul_6_19_g11281/U$1 ( \857 , \824 , \856 );
not \mul_6_19_g11265/U$3 ( \858 , \857 );
xor \mul_6_19_g11418/U$1 ( \859 , \459 , \470 );
xor \mul_6_19_g11418/U$1_r1 ( \860 , \859 , \496 );
not \mul_6_19_g11363/U$3 ( \861 , \860 );
xor \mul_6_19_g11391/U$4 ( \862 , \836 , \838 );
and \mul_6_19_g11391/U$3 ( \863 , \862 , \843 );
and \mul_6_19_g11391/U$5 ( \864 , \836 , \838 );
or \mul_6_19_g11391/U$2 ( \865 , \863 , \864 );
not \mul_6_19_g11390/U$1 ( \866 , \865 );
not \mul_6_19_g11363/U$4 ( \867 , \866 );
or \mul_6_19_g11363/U$2 ( \868 , \861 , \867 );
not \mul_6_19_g11365/U$2 ( \869 , \860 );
nand \mul_6_19_g11365/U$1 ( \870 , \869 , \865 );
nand \mul_6_19_g11363/U$1 ( \871 , \868 , \870 );
xor \mul_6_19_g11375/U$1 ( \872 , \507 , \509 );
xor \mul_6_19_g11375/U$1_r1 ( \873 , \872 , \536 );
xor \g11859/U$1 ( \874 , \871 , \873 );
or \mul_6_19_g11770/U$1 ( \875 , \833 , \829 );
and \mul_6_19_g11349/U$2 ( \876 , \845 , \875 );
and \mul_6_19_g11376/U$2 ( \877 , \829 , \833 );
nor \mul_6_19_g11349/U$1 ( \878 , \876 , \877 );
nand \mul_6_19_g11317/U$1 ( \879 , \874 , \878 );
not \mul_6_19_g11328/U$2 ( \880 , \849 );
not \mul_6_19_g11378/U$1 ( \881 , \853 );
nand \mul_6_19_g11328/U$1 ( \882 , \880 , \881 );
nand \mul_6_19_g11305/U$1 ( \883 , \879 , \882 );
xor \g11878/U$1 ( \884 , \505 , \539 );
xnor \g11878/U$1_r1 ( \885 , \884 , \542 );
not \mul_6_19_g11348/U$3 ( \886 , \860 );
not \mul_6_19_g11348/U$4 ( \887 , \873 );
or \mul_6_19_g11348/U$2 ( \888 , \886 , \887 );
not \mul_6_19_g11389/U$1 ( \889 , \865 );
nand \mul_6_19_g11348/U$1 ( \890 , \888 , \889 );
not \mul_6_19_g11362/U$2 ( \891 , \860 );
not \mul_6_19_g11860/U$1 ( \892 , \873 );
nand \mul_6_19_g11362/U$1 ( \893 , \891 , \892 );
nand \mul_6_19_g11341/U$1 ( \894 , \890 , \893 );
nor \mul_6_19_g11297/U$1 ( \895 , \885 , \894 );
nor \mul_6_19_g11295/U$1 ( \896 , \883 , \895 );
not \mul_6_19_g11265/U$4 ( \897 , \896 );
or \mul_6_19_g11265/U$2 ( \898 , \858 , \897 );
xor \mul_6_19_g11879/U$1 ( \899 , \505 , \539 );
xor \mul_6_19_g11879/U$1_r1 ( \900 , \899 , \542 );
not \mul_6_19_g11335/U$1 ( \901 , \894 );
nand \mul_6_19_g11298/U$1 ( \902 , \900 , \901 );
nor \mul_6_19_g11313/U$1 ( \903 , \874 , \878 );
and \mul_6_19_g11280/U$2 ( \904 , \902 , \903 );
nor \mul_6_19_g11310/U$1 ( \905 , \900 , \901 );
nor \mul_6_19_g11280/U$1 ( \906 , \904 , \905 );
nand \mul_6_19_g11265/U$1 ( \907 , \898 , \906 );
not \mul_6_19_g11249/U$4 ( \908 , \907 );
or \mul_6_19_g11249/U$2 ( \909 , \562 , \908 );
not \mul_6_19_g11279/U$3 ( \910 , \559 );
nor \mul_6_19_g11304/U$1 ( \911 , \503 , \545 );
not \mul_6_19_g11279/U$4 ( \912 , \911 );
or \mul_6_19_g11279/U$2 ( \913 , \910 , \912 );
not \mul_6_19_g11763/U$2 ( \914 , \558 );
nand \mul_6_19_g11763/U$1 ( \915 , \914 , \555 );
nand \mul_6_19_g11279/U$1 ( \916 , \913 , \915 );
nand \mul_6_19_g11268/U$1 ( \917 , \916 , \414 );
not \mul_6_19_g11767/U$2 ( \918 , \412 );
nand \mul_6_19_g11306/U$1 ( \919 , \313 , \357 );
nor \mul_6_19_g11286/U$1 ( \920 , \919 , \386 );
not \mul_6_19_g11766/U$2 ( \921 , \385 );
nor \mul_6_19_g11766/U$1 ( \922 , \921 , \380 );
nor \mul_6_19_g11275/U$1 ( \923 , \920 , \922 );
nor \mul_6_19_g11767/U$1 ( \924 , \918 , \923 );
nor \mul_6_19_g11359/U$1 ( \925 , \409 , \411 );
or \mul_6_19_g11261/U$2 ( \926 , \924 , \925 );
nand \mul_6_19_g11261/U$1 ( \927 , \926 , \405 );
or \mul_6_19_g11398/U$1 ( \928 , \402 , \404 );
and \mul_6_19_g11255/U$1 ( \929 , \917 , \927 , \928 );
nand \mul_6_19_g11249/U$1 ( \930 , \909 , \929 );
not \mul_6_19_g11245/U$4 ( \931 , \930 );
or \mul_6_19_g11245/U$2 ( \932 , \168 , \931 );
or \mul_6_19_g11451/U$1 ( \933 , \165 , \166 );
nand \mul_6_19_g11245/U$1 ( \934 , \932 , \933 );
nand \mul_6_19_g11431/U$1 ( \935 , \167 , \933 );
not \mul_6_19_g11246/U$3 ( \936 , \935 );
not \mul_6_19_g11246/U$4 ( \937 , \930 );
or \mul_6_19_g11246/U$2 ( \938 , \936 , \937 );
or \mul_6_19_g11246/U$5 ( \939 , \935 , \930 );
nand \mul_6_19_g11246/U$1 ( \940 , \938 , \939 );
not \mul_6_19_g11250/U$3 ( \941 , \412 );
nor \mul_6_19_g11272/U$1 ( \942 , \560 , \388 );
not \mul_6_19_g11258/U$3 ( \943 , \942 );
not \mul_6_19_g11258/U$4 ( \944 , \907 );
or \mul_6_19_g11258/U$2 ( \945 , \943 , \944 );
and \g11857/U$1 ( \946 , \358 , \387 );
and \mul_6_19_g11264/U$2 ( \947 , \916 , \946 );
not \mul_6_19_g11274/U$1 ( \948 , \923 );
nor \mul_6_19_g11264/U$1 ( \949 , \947 , \948 );
nand \mul_6_19_g11258/U$1 ( \950 , \945 , \949 );
not \mul_6_19_g11250/U$4 ( \951 , \950 );
or \mul_6_19_g11250/U$2 ( \952 , \941 , \951 );
not \mul_6_19_g11358/U$1 ( \953 , \925 );
nand \mul_6_19_g11250/U$1 ( \954 , \952 , \953 );
nand \mul_6_19_g11384/U$1 ( \955 , \405 , \928 );
not \mul_6_19_g11383/U$1 ( \956 , \955 );
and \mul_6_19_g11247/U$2 ( \957 , \954 , \956 );
not \mul_6_19_g11247/U$4 ( \958 , \954 );
and \mul_6_19_g11247/U$3 ( \959 , \958 , \955 );
nor \mul_6_19_g11247/U$1 ( \960 , \957 , \959 );
buf \fopt11922/U$1 ( \961 , \358 );
not \mul_6_19_g11251/U$3 ( \962 , \961 );
not \mul_6_19_g11293/U$1 ( \963 , \560 );
not \mul_6_19_g11257/U$3 ( \964 , \963 );
not \mul_6_19_g11257/U$4 ( \965 , \907 );
or \mul_6_19_g11257/U$2 ( \966 , \964 , \965 );
not \fopt/U$1 ( \967 , \916 );
nand \mul_6_19_g11257/U$1 ( \968 , \966 , \967 );
not \mul_6_19_g11251/U$4 ( \969 , \968 );
or \mul_6_19_g11251/U$2 ( \970 , \962 , \969 );
buf \fopt11892/U$1 ( \971 , \919 );
nand \mul_6_19_g11251/U$1 ( \972 , \970 , \971 );
not \g11950/U$2 ( \973 , \387 );
nor \g11950/U$1 ( \974 , \973 , \922 );
and \mul_6_19_g11248/U$2 ( \975 , \972 , \974 );
not \mul_6_19_g11248/U$4 ( \976 , \972 );
not \mul_6_19_g11329/U$1 ( \977 , \974 );
and \mul_6_19_g11248/U$3 ( \978 , \976 , \977 );
nor \mul_6_19_g11248/U$1 ( \979 , \975 , \978 );
buf \fopt11921/U$1 ( \980 , \546 );
not \mul_6_19_g11259/U$3 ( \981 , \980 );
not \mul_6_19_g11259/U$4 ( \982 , \907 );
or \mul_6_19_g11259/U$2 ( \983 , \981 , \982 );
not \mul_6_19_g11303/U$1 ( \984 , \911 );
nand \mul_6_19_g11259/U$1 ( \985 , \983 , \984 );
nand \mul_6_19_g11289/U$1 ( \986 , \559 , \915 );
not \mul_6_19_g11288/U$1 ( \987 , \986 );
and \mul_6_19_g11254/U$2 ( \988 , \985 , \987 );
not \mul_6_19_g11254/U$4 ( \989 , \985 );
and \mul_6_19_g11254/U$3 ( \990 , \989 , \986 );
nor \mul_6_19_g11254/U$1 ( \991 , \988 , \990 );
nand \mul_6_19_g11270/U$1 ( \992 , \857 , \882 );
not \mul_6_19_g11269/U$1 ( \993 , \992 );
buf \mul_6_19_g11316/U$1 ( \994 , \879 );
and \mul_6_19_g11262/U$2 ( \995 , \993 , \994 );
buf \fopt11900/U$1 ( \996 , \903 );
nor \mul_6_19_g11262/U$1 ( \997 , \995 , \996 );
not \mul_6_19_g11292/U$2 ( \998 , \905 );
nand \mul_6_19_g11292/U$1 ( \999 , \998 , \902 );
and \mul_6_19_g11256/U$2 ( \1000 , \997 , \999 );
not \mul_6_19_g11256/U$4 ( \1001 , \997 );
not \mul_6_19_g11291/U$1 ( \1002 , \999 );
and \mul_6_19_g11256/U$3 ( \1003 , \1001 , \1002 );
nor \mul_6_19_g11256/U$1 ( \1004 , \1000 , \1003 );
not \fopt11899/U$1 ( \1005 , \996 );
nand \mul_6_19_g11308/U$1 ( \1006 , \1005 , \994 );
and \mul_6_19_g11263/U$2 ( \1007 , \992 , \1006 );
not \mul_6_19_g11263/U$4 ( \1008 , \992 );
not \mul_6_19_g11307/U$1 ( \1009 , \1006 );
and \mul_6_19_g11263/U$3 ( \1010 , \1008 , \1009 );
nor \mul_6_19_g11263/U$1 ( \1011 , \1007 , \1010 );
nand \mul_6_19_g11273/U$1 ( \1012 , \824 , \855 );
nand \mul_6_19_g11319/U$1 ( \1013 , \882 , \854 );
not \mul_6_19_g11318/U$1 ( \1014 , \1013 );
and \mul_6_19_g11266/U$2 ( \1015 , \1012 , \1014 );
not \mul_6_19_g11266/U$4 ( \1016 , \1012 );
and \mul_6_19_g11266/U$3 ( \1017 , \1016 , \1013 );
nor \mul_6_19_g11266/U$1 ( \1018 , \1015 , \1017 );
nand \mul_6_19_g11346/U$1 ( \1019 , \823 , \855 );
not \mul_6_19_g11345/U$1 ( \1020 , \1019 );
and \mul_6_19_g11282/U$2 ( \1021 , \770 , \1020 );
not \mul_6_19_g11282/U$4 ( \1022 , \770 );
and \mul_6_19_g11282/U$3 ( \1023 , \1022 , \1019 );
nor \mul_6_19_g11282/U$1 ( \1024 , \1021 , \1023 );
nand \mul_6_19_g11287/U$1 ( \1025 , \961 , \971 );
nand \mul_6_19_g11290/U$1 ( \1026 , \984 , \980 );
nand \mul_6_19_g11368/U$1 ( \1027 , \769 , \665 );
not \mul_6_19_g11321/U$3 ( \1028 , \1027 );
buf \mul_6_19_g11342/U$1 ( \1029 , \764 );
not \mul_6_19_g11321/U$4 ( \1030 , \1029 );
or \mul_6_19_g11321/U$2 ( \1031 , \1028 , \1030 );
or \mul_6_19_g11321/U$5 ( \1032 , \1029 , \1027 );
nand \mul_6_19_g11321/U$1 ( \1033 , \1031 , \1032 );
nand \mul_6_19_g11347/U$1 ( \1034 , \412 , \953 );
buf \mul_6_19_g11369/U$1 ( \1035 , \758 );
not \mul_6_19_g11352/U$3 ( \1036 , \1035 );
nand \mul_6_19_g11382/U$1 ( \1037 , \763 , \684 );
not \mul_6_19_g11352/U$4 ( \1038 , \1037 );
or \mul_6_19_g11352/U$2 ( \1039 , \1036 , \1038 );
or \mul_6_19_g11352/U$5 ( \1040 , \1035 , \1037 );
nand \mul_6_19_g11352/U$1 ( \1041 , \1039 , \1040 );
and \mul_6_19_g11771/U$1 ( \1042 , \757 , \703 );
and \mul_6_19_g11386/U$2 ( \1043 , \1042 , \754 );
not \mul_6_19_g11386/U$4 ( \1044 , \1042 );
not \mul_6_19_g11406/U$1 ( \1045 , \754 );
and \mul_6_19_g11386/U$3 ( \1046 , \1044 , \1045 );
nor \mul_6_19_g11386/U$1 ( \1047 , \1043 , \1046 );
nand \mul_6_19_g11432/U$1 ( \1048 , \721 , \752 );
not \mul_6_19_g11437/U$1 ( \1049 , \751 );
and \mul_6_19_g11417/U$2 ( \1050 , \1048 , \1049 );
not \mul_6_19_g11417/U$4 ( \1051 , \1048 );
and \mul_6_19_g11417/U$3 ( \1052 , \1051 , \751 );
nor \mul_6_19_g11417/U$1 ( \1053 , \1050 , \1052 );
nand \mul_6_19_g11483/U$1 ( \1054 , \750 , \736 );
not \mul_6_19_g11460/U$3 ( \1055 , \1054 );
not \mul_6_19_g11460/U$4 ( \1056 , \746 );
or \mul_6_19_g11460/U$2 ( \1057 , \1055 , \1056 );
or \mul_6_19_g11460/U$5 ( \1058 , \746 , \1054 );
nand \mul_6_19_g11460/U$1 ( \1059 , \1057 , \1058 );
xor \mul_6_19_g11484/U$1 ( \1060 , \739 , \741 );
xor \mul_6_19_g11484/U$1_r1 ( \1061 , \1060 , \743 );
and \mul_6_19_g11618/U$2 ( \1062 , \111 , \B[0] );
and \mul_6_19_g11618/U$3 ( \1063 , \118 , \B[1] );
nor \mul_6_19_g11618/U$1 ( \1064 , \1062 , \1063 );
nor \mul_6_19_g11579/U$1 ( \1065 , \741 , \1064 );
not \mul_6_19_g11644/U$1 ( \1066 , \740 );
xnor \g2/U$1 ( \1067 , \950 , \1034 );
xnor \g11791/U$1 ( \1068 , \968 , \1025 );
xnor \g11792/U$1 ( \1069 , \1026 , \907 );
endmodule

